///////////////////////////////////////////////////////////////////////////////
//  Copyright 2018 Fredrik A. Kristiansen
//  Permission is hereby granted, free of charge, to any person obtaining a 
//  copy of this software and associated documentation files (the "Software"), 
//  to deal in the Software without restriction, including without limitation 
//  the rights to use, copy, modify, merge, publish, distribute, sublicense, 
//  and/or sell copies of the Software, and to permit persons to whom the 
//  Software is furnished to do so, subject to the following conditions:
//
//  The above copyright notice and this permission notice shall be included in 
//  all copies or substantial portions of the Software.
//
//  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS 
//  OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
//  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE 
//  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER 
//  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
//  FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER 
//  DEALINGS IN THE SOFTWARE.
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps
`include "interrupt_encoder.v"

module interrupt_encoder_tb();
	reg  [6:0] irq_n;
	wire [2:0] ipl_n;

	interrupt_encoder encoder(
		.a_n(irq_n),
		.y_n(ipl_n)
	);

	initial begin
		$dumpfile("interrupt_encoder_tb.vcd");
		$dumpvars(0, encoder);

		irq_n = 7'b1111111;
		#1 irq_n = 7'b0101011;
		#1 irq_n = 7'b0111111;
		#1 irq_n = 7'b1110101;
		#1 irq_n = 7'b1111110;
		#1 $finish;
	end
endmodule
